.include subs.cir
*lcon is very important.
.param Lcon=.1p
.param Vmag=0.95* 548m
*1.1 works
.param Vfreq=1G
*V = phi0/ (C 2pi f 2L) = 2.067E-15 / (10^-13 6.28)
.param Imag=1m
.param shift=166p
*Imag -.6 w L = 1.46
* clock network meanders

*Vex0       1    0     sin(0 Vmag Vfreq)
*Vex90      2    0     sin(0 Vmag Vfreq shift)
*Vex180     3    0     sin(0 Vmag Vfreq 2*shift)
*Vex270     4    0     sin(0 Vmag Vfreq 3*shift)

* alternate network
*seems 8 phases is necessary.
*the hypothesis is that this is because a junction switches with the absolute magnitude of the clock current, which comes around with double the frequency of the clock.
*This means we need 4 networks, both with positive and negative leads.

*Iex1       21    22     sin(0 Imag Vfreq)
*Iex2       23    24     sin(0 Imag Vfreq shift)
*Iex3       25    26     sin(0 Imag Vfreq 2*shift)
*Iex4       27    28     sin(0 Imag Vfreq 3*shift)
*Iex5       29    30     sin(0 Imag Vfreq 4*shift)

*C1 C2 Lin Louts
*X1 cbuf 21 22 5 6 
*X2 cbuf 23 24 7 8
*X3 cbuf 25 26 9 10
*X4 cbuf 27 28 11 12
*X5 cbuf 29 30 13 14

  
*another test clock.
*only 3*2 clocks are needed it seems.

V0       31    0     sin(0 Vmag Vfreq 0)
V_60     32    0     sin(0 Vmag Vfreq -5*shift)
V_120    33    0     sin(0 Vmag Vfreq -4*shift)
V_180    34    0     sin(0 Vmag Vfreq -3*shift)
V_240    35    0     sin(0 Vmag Vfreq -2*shift)
V_300    36    0     sin(0 Vmag Vfreq -1*shift)


X1 cbuf 31 34 5 6 
X2 cbuf 32 35 7 8
X3 cbuf 33 36 9 10
X4 cbuf 34 31 11 12
X5 cbuf 35 32 13 14
x6 cbuf 36 33 15 16

X7 cbuf 31 34 17 18
X8 cbuf 32 35 19 20
X9 cbuf 33 36 21 22
X10 cbuf 34 31 23 24
X11 cbuf 35 32 25 26
x12 cbuf 36 33 27 28

*Iin1       0    5      pwl(0 10u .95n 10u 1.05n -10u 2n -10u)
*Iin1       0    5      10u
*Iin1       0    5       pwl(0 -20u 2.99n -20u 3n 20u 3.99n 20u 4n -20u)
Iin       0    5       cus(wform.txt .25p 1u)


Lcon1   6   7   Lcon
Lcon2   8   9   Lcon       
Lcon3   10  11  Lcon
Lcon4   12  13  Lcon
Lcon5   14  15  Lcon

Lcon6   16  17   Lcon
Lcon7   18  19   Lcon       
Lcon8   20  21  Lcon
Lcon9   22  23  Lcon
Lcon10  24  25  Lcon
Lcon11  26  27  Lcon
Lout    28  0   20p

.tran .25p 12n 1n 11p


.print DEVI V0
.print DEVI Iin

*.print DEVV Vex0
*.print DEVI B1.X3
*.print DEVV B1.X3
.print DEVI Lst.X1
*.print DEVI Lcon1
*.print DEVI Lst.X2
*.print DEVI Lcon2
*.print DEVI Lst.X3
*.print DEVI Lcon3
*.print DEVI Lst.X4
*.print DEVI Lcon4
.print DEVI Lst.X5
*.print DEVI Lcon5
.print DEVI Lst.X6
*.print DEVI Lst.X7
*.print DEVI Lst.X8
*.print DEVI Lst.X9
*.print DEVI Lst.X10
*.print DEVI Lst.X11
.print DEVI Lst.X12
*.print DEVI Lcon2
*.print DEVI Lcon3
*.print DEVI Lcon4
.print DEVI Lout

.end