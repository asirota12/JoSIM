.include subs.cir
*lcon is very important.
.param Lcon=.1p
.param Vmag=500m
*1000m with 1.46 L
.param Vfreq=1G
.param Imag=.4m
.param shift=166p
*Imag -.6 w L = 1.46

* I would like to make a plot of the output current vs the through current


* clock network meanders

Icross1    31    0    pwl(0 0 1n 0 3n Imag)
Icross2    34    0    pwl(0 0 1n 0 3n -Imag)

*Pcross1    31    0    pwl(0 0 1n 0 3n Imag)
*Pcross2    34    0    pwl(0 0 1n 0 3n -Imag)


X1 cbuf 31 34 1 2 

*Iin1       0    5      pwl(0 10u .95n 10u 1.05n -10u 2n -10u)
*Iin1       0    5      10u
*Iin1       0    5       pwl(0 -20u 2.99n -20u 3n 20u 3.99n 20u 4n -20u)
Iin1       0    1       cus(wform.txt .25p 1u)

Lout    2  0   .1p

.tran .25p 3n 1n 10p

*.print DEVI Iex1
*.print DEVI Iex2

.print DEVI Icross1
.print DEVI Iin1

.print DEVI Lst.X1
.print DEVI L1.X1
.print DEVI LG1.X1
.print DEVI L2.X1
.print DEVI LG2.X1
.print NODEP 3.X1
.print NODEP 5.X1
*.print DEVI Lout

.end
